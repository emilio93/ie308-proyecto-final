**************************************
*      DIODO ZENER 1N4733            *
**************************************
.MODEL 1n4733 d(
  + BV=5.1
  + IBV=49m
  + Rs=7
  + Is=1.214f
  + Ikf=0
  + N=1
  + Xti=3
  + Eg=1.1
  + Cjo=185p
  + M=.3509
  + Vj=.75
  + Fc=.5
  + Nbv=.74348)
