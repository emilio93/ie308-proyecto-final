*
.SUBCKT LM317 1 2 3
  * IN OUT ADJ
  IADJ 1 4 50U
  VREF 4 3 1.25
  RC 1 14 0.742
  DBK 14 13 D1
  CBC 13 15 2.479N
  RBC 15 5 247
  QP 13 5 2 Q1
  RB2 6 5 124
  DSC 6 11 D1
  ESC 11 2 POLY(2) (13,5) (6,5) 2.85
  + 0 0 0 -70.1M
  DFB 6 12 D1
  EFB 12 2 POLY(2) (13,5) (6,5) 3.92
  + -135M 0 1.21M -70.1M
  RB1 7 6 1
  EB 7 2 8 2 2.56
  CPZ 10 2 0.796U
  DPU 10 2 D1
  RZ 8 10 0.104
  RP 9 8 100
  EP 9 2 4 2 103.6
  RI 2 4 100MEG
  .MODEL Q1 NPN (IS=30F BF=100
  + VAF=14.27 NF=1.604)
  .MODEL D1 D (IS=30F N=1.604)
.ENDS LM317
