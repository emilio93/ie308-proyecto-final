
.SUBCKT LM337K 8 1 19
*Connections Input Adj. Output
*LM337 negative voltage regulator
.MODEL QN NPN (BF=50 TF=1N CJC=1P)
.MODEL QPOUT PNP (BF=50 TF=1N RE=.2 CJC=1P)
.MODEL QP PNP CJC=1P TF=2N
.MODEL DN D
.MODEL D2 D BV=12 IBV=100U
R10 25 6 1K
Q3 8 17 16 QPOUT
Q4 8 25 17 QP
R18 19 17 250
R19 19 16 .3
G1 8 6 1 18 .1
C7 6 2 .04U
R24 2 8 100
I_ADJ 0 1 65U
R26 8 25 200K
Q5 25 4 19 QP
R27 16 4 200
R28 7 4 7K
D1 8 7 D2
D2 8 6 DN
V1 18 19 1.25
.ENDS
************
